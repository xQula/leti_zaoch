library verilog;
use verilog.vl_types.all;
entity jk_trig_vlg_vec_tst is
end jk_trig_vlg_vec_tst;
