library verilog;
use verilog.vl_types.all;
entity d_trig_vlg_vec_tst is
end d_trig_vlg_vec_tst;
