library verilog;
use verilog.vl_types.all;
entity lab_4_multireg_vlg_vec_tst is
end lab_4_multireg_vlg_vec_tst;
