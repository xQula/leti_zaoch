library verilog;
use verilog.vl_types.all;
entity t_trig_vlg_vec_tst is
end t_trig_vlg_vec_tst;
